`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: and
// Description: 2-input AND gate
//////////////////////////////////////////////////////////////////////////////////

module and_gate (
    input A,
    input B,
    output C
);

    assign C = A & B;

endmodule
